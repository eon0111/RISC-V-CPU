module ALU(
  input  [3:0]  io_func, // @[ca2023-lab3/src/main/scala/riscv/core/ALU.scala 16:14]
  input  [31:0] io_op1, // @[ca2023-lab3/src/main/scala/riscv/core/ALU.scala 16:14]
  input  [31:0] io_op2, // @[ca2023-lab3/src/main/scala/riscv/core/ALU.scala 16:14]
  output [31:0] io_result // @[ca2023-lab3/src/main/scala/riscv/core/ALU.scala 16:14]
);
  wire [31:0] _io_result_T_1 = io_op1 + io_op2; // @[ca2023-lab3/src/main/scala/riscv/core/ALU.scala 28:27]
  wire [31:0] _io_result_T_3 = io_op1 - io_op2; // @[ca2023-lab3/src/main/scala/riscv/core/ALU.scala 31:27]
  wire [62:0] _GEN_10 = {{31'd0}, io_op1}; // @[ca2023-lab3/src/main/scala/riscv/core/ALU.scala 34:27]
  wire [62:0] _io_result_T_5 = _GEN_10 << io_op2[4:0]; // @[ca2023-lab3/src/main/scala/riscv/core/ALU.scala 34:27]
  wire [31:0] _io_result_T_6 = io_op1; // @[ca2023-lab3/src/main/scala/riscv/core/ALU.scala 37:27]
  wire [31:0] _io_result_T_7 = io_op2; // @[ca2023-lab3/src/main/scala/riscv/core/ALU.scala 37:43]
  wire [31:0] _io_result_T_9 = io_op1 ^ io_op2; // @[ca2023-lab3/src/main/scala/riscv/core/ALU.scala 40:27]
  wire [31:0] _io_result_T_10 = io_op1 | io_op2; // @[ca2023-lab3/src/main/scala/riscv/core/ALU.scala 43:27]
  wire [31:0] _io_result_T_11 = io_op1 & io_op2; // @[ca2023-lab3/src/main/scala/riscv/core/ALU.scala 46:27]
  wire [31:0] _io_result_T_13 = io_op1 >> io_op2[4:0]; // @[ca2023-lab3/src/main/scala/riscv/core/ALU.scala 49:27]
  wire [31:0] _io_result_T_17 = $signed(io_op1) >>> io_op2[4:0]; // @[ca2023-lab3/src/main/scala/riscv/core/ALU.scala 52:52]
  wire  _GEN_0 = 4'ha == io_func & io_op1 < io_op2; // @[ca2023-lab3/src/main/scala/riscv/core/ALU.scala 25:13 26:19 55:17]
  wire [31:0] _GEN_1 = 4'h9 == io_func ? _io_result_T_17 : {{31'd0}, _GEN_0}; // @[ca2023-lab3/src/main/scala/riscv/core/ALU.scala 26:19 52:17]
  wire [31:0] _GEN_2 = 4'h8 == io_func ? _io_result_T_13 : _GEN_1; // @[ca2023-lab3/src/main/scala/riscv/core/ALU.scala 26:19 49:17]
  wire [31:0] _GEN_3 = 4'h7 == io_func ? _io_result_T_11 : _GEN_2; // @[ca2023-lab3/src/main/scala/riscv/core/ALU.scala 26:19 46:17]
  wire [31:0] _GEN_4 = 4'h6 == io_func ? _io_result_T_10 : _GEN_3; // @[ca2023-lab3/src/main/scala/riscv/core/ALU.scala 26:19 43:17]
  wire [31:0] _GEN_5 = 4'h5 == io_func ? _io_result_T_9 : _GEN_4; // @[ca2023-lab3/src/main/scala/riscv/core/ALU.scala 26:19 40:17]
  wire [31:0] _GEN_6 = 4'h4 == io_func ? {{31'd0}, $signed(_io_result_T_6) < $signed(_io_result_T_7)} : _GEN_5; // @[ca2023-lab3/src/main/scala/riscv/core/ALU.scala 26:19 37:17]
  wire [62:0] _GEN_7 = 4'h3 == io_func ? _io_result_T_5 : {{31'd0}, _GEN_6}; // @[ca2023-lab3/src/main/scala/riscv/core/ALU.scala 26:19 34:17]
  wire [62:0] _GEN_8 = 4'h2 == io_func ? {{31'd0}, _io_result_T_3} : _GEN_7; // @[ca2023-lab3/src/main/scala/riscv/core/ALU.scala 26:19 31:17]
  wire [62:0] _GEN_9 = 4'h1 == io_func ? {{31'd0}, _io_result_T_1} : _GEN_8; // @[ca2023-lab3/src/main/scala/riscv/core/ALU.scala 26:19 28:17]
  assign io_result = _GEN_9[31:0];
endmodule
module ALUControl(
  input  [6:0] io_opcode, // @[ca2023-lab3/src/main/scala/riscv/core/ALUControl.scala 10:14]
  input  [2:0] io_funct3, // @[ca2023-lab3/src/main/scala/riscv/core/ALUControl.scala 10:14]
  input  [6:0] io_funct7, // @[ca2023-lab3/src/main/scala/riscv/core/ALUControl.scala 10:14]
  output [3:0] io_alu_funct // @[ca2023-lab3/src/main/scala/riscv/core/ALUControl.scala 10:14]
);
  wire [3:0] _io_alu_funct_T_1 = io_funct7[5] ? 4'h9 : 4'h8; // @[ca2023-lab3/src/main/scala/riscv/core/ALUControl.scala 33:41]
  wire [1:0] _io_alu_funct_T_3 = 3'h1 == io_funct3 ? 2'h3 : 2'h1; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire [2:0] _io_alu_funct_T_5 = 3'h2 == io_funct3 ? 3'h4 : {{1'd0}, _io_alu_funct_T_3}; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire [3:0] _io_alu_funct_T_7 = 3'h3 == io_funct3 ? 4'ha : {{1'd0}, _io_alu_funct_T_5}; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire [3:0] _io_alu_funct_T_9 = 3'h4 == io_funct3 ? 4'h5 : _io_alu_funct_T_7; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire [3:0] _io_alu_funct_T_11 = 3'h6 == io_funct3 ? 4'h6 : _io_alu_funct_T_9; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire [3:0] _io_alu_funct_T_13 = 3'h7 == io_funct3 ? 4'h7 : _io_alu_funct_T_11; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire [3:0] _io_alu_funct_T_15 = 3'h5 == io_funct3 ? _io_alu_funct_T_1 : _io_alu_funct_T_13; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire [1:0] _io_alu_funct_T_17 = io_funct7[5] ? 2'h2 : 2'h1; // @[ca2023-lab3/src/main/scala/riscv/core/ALUControl.scala 42:43]
  wire [1:0] _io_alu_funct_T_21 = 3'h1 == io_funct3 ? 2'h3 : _io_alu_funct_T_17; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire [2:0] _io_alu_funct_T_23 = 3'h2 == io_funct3 ? 3'h4 : {{1'd0}, _io_alu_funct_T_21}; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire [3:0] _io_alu_funct_T_25 = 3'h3 == io_funct3 ? 4'ha : {{1'd0}, _io_alu_funct_T_23}; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire [3:0] _io_alu_funct_T_27 = 3'h4 == io_funct3 ? 4'h5 : _io_alu_funct_T_25; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire [3:0] _io_alu_funct_T_29 = 3'h6 == io_funct3 ? 4'h6 : _io_alu_funct_T_27; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire [3:0] _io_alu_funct_T_31 = 3'h7 == io_funct3 ? 4'h7 : _io_alu_funct_T_29; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire [3:0] _io_alu_funct_T_33 = 3'h5 == io_funct3 ? _io_alu_funct_T_1 : _io_alu_funct_T_31; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _GEN_1 = 7'h37 == io_opcode | 7'h17 == io_opcode; // @[ca2023-lab3/src/main/scala/riscv/core/ALUControl.scala 20:21 69:20]
  wire  _GEN_2 = 7'h67 == io_opcode | _GEN_1; // @[ca2023-lab3/src/main/scala/riscv/core/ALUControl.scala 20:21 66:20]
  wire  _GEN_3 = 7'h6f == io_opcode | _GEN_2; // @[ca2023-lab3/src/main/scala/riscv/core/ALUControl.scala 20:21 63:20]
  wire  _GEN_4 = 7'h23 == io_opcode | _GEN_3; // @[ca2023-lab3/src/main/scala/riscv/core/ALUControl.scala 20:21 60:20]
  wire  _GEN_5 = 7'h3 == io_opcode | _GEN_4; // @[ca2023-lab3/src/main/scala/riscv/core/ALUControl.scala 20:21 57:20]
  wire  _GEN_6 = 7'h63 == io_opcode | _GEN_5; // @[ca2023-lab3/src/main/scala/riscv/core/ALUControl.scala 20:21 54:20]
  wire [3:0] _GEN_7 = 7'h33 == io_opcode ? _io_alu_funct_T_33 : {{3'd0}, _GEN_6}; // @[ca2023-lab3/src/main/scala/riscv/core/ALUControl.scala 20:21 38:20]
  assign io_alu_funct = 7'h13 == io_opcode ? _io_alu_funct_T_15 : _GEN_7; // @[ca2023-lab3/src/main/scala/riscv/core/ALUControl.scala 20:21 22:20]
endmodule
module Execute(
  input         clock,
  input         reset,
  input  [31:0] io_instruction, // @[home/eon/Documentos/TFM/RISC-V-CPU/ca2023-lab3/src/main/scala/riscv/core/Execute.scala 13:14]
  input  [31:0] io_instruction_address, // @[home/eon/Documentos/TFM/RISC-V-CPU/ca2023-lab3/src/main/scala/riscv/core/Execute.scala 13:14]
  input  [31:0] io_reg1_data, // @[home/eon/Documentos/TFM/RISC-V-CPU/ca2023-lab3/src/main/scala/riscv/core/Execute.scala 13:14]
  input  [31:0] io_reg2_data, // @[home/eon/Documentos/TFM/RISC-V-CPU/ca2023-lab3/src/main/scala/riscv/core/Execute.scala 13:14]
  input  [31:0] io_immediate, // @[home/eon/Documentos/TFM/RISC-V-CPU/ca2023-lab3/src/main/scala/riscv/core/Execute.scala 13:14]
  input         io_aluop1_source, // @[home/eon/Documentos/TFM/RISC-V-CPU/ca2023-lab3/src/main/scala/riscv/core/Execute.scala 13:14]
  input         io_aluop2_source, // @[home/eon/Documentos/TFM/RISC-V-CPU/ca2023-lab3/src/main/scala/riscv/core/Execute.scala 13:14]
  output [31:0] io_mem_alu_result, // @[home/eon/Documentos/TFM/RISC-V-CPU/ca2023-lab3/src/main/scala/riscv/core/Execute.scala 13:14]
  output        io_if_jump_flag, // @[home/eon/Documentos/TFM/RISC-V-CPU/ca2023-lab3/src/main/scala/riscv/core/Execute.scala 13:14]
  output [31:0] io_if_jump_address // @[home/eon/Documentos/TFM/RISC-V-CPU/ca2023-lab3/src/main/scala/riscv/core/Execute.scala 13:14]
);
  wire [3:0] alu_io_func; // @[home/eon/Documentos/TFM/RISC-V-CPU/ca2023-lab3/src/main/scala/riscv/core/Execute.scala 33:24]
  wire [31:0] alu_io_op1; // @[home/eon/Documentos/TFM/RISC-V-CPU/ca2023-lab3/src/main/scala/riscv/core/Execute.scala 33:24]
  wire [31:0] alu_io_op2; // @[home/eon/Documentos/TFM/RISC-V-CPU/ca2023-lab3/src/main/scala/riscv/core/Execute.scala 33:24]
  wire [31:0] alu_io_result; // @[home/eon/Documentos/TFM/RISC-V-CPU/ca2023-lab3/src/main/scala/riscv/core/Execute.scala 33:24]
  wire [6:0] alu_ctrl_io_opcode; // @[home/eon/Documentos/TFM/RISC-V-CPU/ca2023-lab3/src/main/scala/riscv/core/Execute.scala 34:24]
  wire [2:0] alu_ctrl_io_funct3; // @[home/eon/Documentos/TFM/RISC-V-CPU/ca2023-lab3/src/main/scala/riscv/core/Execute.scala 34:24]
  wire [6:0] alu_ctrl_io_funct7; // @[home/eon/Documentos/TFM/RISC-V-CPU/ca2023-lab3/src/main/scala/riscv/core/Execute.scala 34:24]
  wire [3:0] alu_ctrl_io_alu_funct; // @[home/eon/Documentos/TFM/RISC-V-CPU/ca2023-lab3/src/main/scala/riscv/core/Execute.scala 34:24]
  wire [6:0] opcode = io_instruction[6:0]; // @[home/eon/Documentos/TFM/RISC-V-CPU/ca2023-lab3/src/main/scala/riscv/core/Execute.scala 27:30]
  wire [2:0] funct3 = io_instruction[14:12]; // @[home/eon/Documentos/TFM/RISC-V-CPU/ca2023-lab3/src/main/scala/riscv/core/Execute.scala 28:30]
  wire  _io_if_jump_flag_T_1 = opcode == 7'h67; // @[home/eon/Documentos/TFM/RISC-V-CPU/ca2023-lab3/src/main/scala/riscv/core/Execute.scala 61:13]
  wire  _io_if_jump_flag_T_2 = opcode == 7'h6f | _io_if_jump_flag_T_1; // @[home/eon/Documentos/TFM/RISC-V-CPU/ca2023-lab3/src/main/scala/riscv/core/Execute.scala 60:50]
  wire  _io_if_jump_flag_T_4 = io_reg1_data == io_reg2_data; // @[home/eon/Documentos/TFM/RISC-V-CPU/ca2023-lab3/src/main/scala/riscv/core/Execute.scala 66:49]
  wire  _io_if_jump_flag_T_5 = io_reg1_data != io_reg2_data; // @[home/eon/Documentos/TFM/RISC-V-CPU/ca2023-lab3/src/main/scala/riscv/core/Execute.scala 67:49]
  wire  _io_if_jump_flag_T_8 = $signed(io_reg1_data) < $signed(io_reg2_data); // @[home/eon/Documentos/TFM/RISC-V-CPU/ca2023-lab3/src/main/scala/riscv/core/Execute.scala 68:56]
  wire  _io_if_jump_flag_T_11 = $signed(io_reg1_data) >= $signed(io_reg2_data); // @[home/eon/Documentos/TFM/RISC-V-CPU/ca2023-lab3/src/main/scala/riscv/core/Execute.scala 69:56]
  wire  _io_if_jump_flag_T_12 = io_reg1_data < io_reg2_data; // @[home/eon/Documentos/TFM/RISC-V-CPU/ca2023-lab3/src/main/scala/riscv/core/Execute.scala 70:56]
  wire  _io_if_jump_flag_T_13 = io_reg1_data >= io_reg2_data; // @[home/eon/Documentos/TFM/RISC-V-CPU/ca2023-lab3/src/main/scala/riscv/core/Execute.scala 71:56]
  wire  _io_if_jump_flag_T_17 = 3'h1 == funct3 ? _io_if_jump_flag_T_5 : 3'h0 == funct3 & _io_if_jump_flag_T_4; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _io_if_jump_flag_T_19 = 3'h4 == funct3 ? _io_if_jump_flag_T_8 : _io_if_jump_flag_T_17; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _io_if_jump_flag_T_21 = 3'h5 == funct3 ? _io_if_jump_flag_T_11 : _io_if_jump_flag_T_19; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _io_if_jump_flag_T_23 = 3'h6 == funct3 ? _io_if_jump_flag_T_12 : _io_if_jump_flag_T_21; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _io_if_jump_flag_T_25 = 3'h7 == funct3 ? _io_if_jump_flag_T_13 : _io_if_jump_flag_T_23; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _io_if_jump_flag_T_26 = opcode == 7'h63 & _io_if_jump_flag_T_25; // @[home/eon/Documentos/TFM/RISC-V-CPU/ca2023-lab3/src/main/scala/riscv/core/Execute.scala 62:37]
  wire [31:0] _io_if_jump_address_T_1 = _io_if_jump_flag_T_1 ? io_reg1_data : io_instruction_address; // @[home/eon/Documentos/TFM/RISC-V-CPU/ca2023-lab3/src/main/scala/riscv/core/Execute.scala 74:43]
  ALU alu ( // @[home/eon/Documentos/TFM/RISC-V-CPU/ca2023-lab3/src/main/scala/riscv/core/Execute.scala 33:24]
    .io_func(alu_io_func),
    .io_op1(alu_io_op1),
    .io_op2(alu_io_op2),
    .io_result(alu_io_result)
  );
  ALUControl alu_ctrl ( // @[home/eon/Documentos/TFM/RISC-V-CPU/ca2023-lab3/src/main/scala/riscv/core/Execute.scala 34:24]
    .io_opcode(alu_ctrl_io_opcode),
    .io_funct3(alu_ctrl_io_funct3),
    .io_funct7(alu_ctrl_io_funct7),
    .io_alu_funct(alu_ctrl_io_alu_funct)
  );
  assign io_mem_alu_result = alu_io_result; // @[home/eon/Documentos/TFM/RISC-V-CPU/ca2023-lab3/src/main/scala/riscv/core/Execute.scala 59:21]
  assign io_if_jump_flag = _io_if_jump_flag_T_2 | _io_if_jump_flag_T_26; // @[home/eon/Documentos/TFM/RISC-V-CPU/ca2023-lab3/src/main/scala/riscv/core/Execute.scala 61:36]
  assign io_if_jump_address = io_immediate + _io_if_jump_address_T_1; // @[home/eon/Documentos/TFM/RISC-V-CPU/ca2023-lab3/src/main/scala/riscv/core/Execute.scala 74:38]
  assign alu_io_func = alu_ctrl_io_alu_funct; // @[home/eon/Documentos/TFM/RISC-V-CPU/ca2023-lab3/src/main/scala/riscv/core/Execute.scala 43:15]
  assign alu_io_op1 = io_aluop1_source ? io_instruction_address : io_reg1_data; // @[home/eon/Documentos/TFM/RISC-V-CPU/ca2023-lab3/src/main/scala/riscv/core/Execute.scala 45:20]
  assign alu_io_op2 = io_aluop2_source ? io_immediate : io_reg2_data; // @[home/eon/Documentos/TFM/RISC-V-CPU/ca2023-lab3/src/main/scala/riscv/core/Execute.scala 51:20]
  assign alu_ctrl_io_opcode = io_instruction[6:0]; // @[home/eon/Documentos/TFM/RISC-V-CPU/ca2023-lab3/src/main/scala/riscv/core/Execute.scala 27:30]
  assign alu_ctrl_io_funct3 = io_instruction[14:12]; // @[home/eon/Documentos/TFM/RISC-V-CPU/ca2023-lab3/src/main/scala/riscv/core/Execute.scala 28:30]
  assign alu_ctrl_io_funct7 = io_instruction[31:25]; // @[home/eon/Documentos/TFM/RISC-V-CPU/ca2023-lab3/src/main/scala/riscv/core/Execute.scala 29:30]
endmodule
